module LED_Pixel_Encoder ();
	//TODO: WIP
endmodule // LED_Pixel_Encoder
