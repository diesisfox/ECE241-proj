module Top_Ctrl (
	input CLOCK_50, PS2_CLK, PS2_DAT,
	input [3:0] KEY,
	input [9:0] LEDR,
	input [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5,
	output [1:0] GPIO_0
	);

endmodule // Top_Ctrl
